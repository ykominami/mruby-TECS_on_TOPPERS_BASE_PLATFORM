/*
 *  @(#) $Id: tSerialPort.cdl 439 2009-07-22 09:08:30Z ertl-takuya $
 */

/**** Wrapper ����  *****/
import_C( "syssvc/serial.h" );

/*
 *		���ꥢ�륤�󥿥ե������ɥ饤�ФΥ���ݡ��ͥ�ȵ��ҥե�����
 *
 *      ����� TECS �ǤǤϤʤ�����¸�� ASP �� serial ��ñ��ʥ�åѡ��Ǥ��롥
 *      ��ü���᤯ tSample ��¸����뤿��ˡ���åѡ��Ȥ��Ƥ��롥
 */

// +-----------------------------
// typedef struct {
// 	uint_t		reacnt;				/* �����Хåե����ʸ���� */
// 	uint_t		wricnt;				/* �����Хåե����ʸ���� */
// } T_SERIAL_RPOR;
// -----------------------------+

signature sSerialPort {
	ER		open(void);
	ER		close(void);
	ER_UINT	read([out,size_is(length)] char_t *buffer, [in] uint_t length);
	ER_UINT	write([in,size_is(length)] const char_t *buffer, [in] uint_t length);
	ER		control([in] uint_t ioControl);
	ER		refer([out] T_SERIAL_RPOR *pk_rpor);
};

signature snSerialPort {
	bool_t	getChar([out] char_t *p_char);
};

// +------------------------------------------
// /* ���ꥢ�륤�󥿥ե������ɥ饤�Ф�ư�������ѤΤ������� */
// const uint_t IOCTL_NULL	= 0;		/* ����ʤ� */
// const uint_t IOCTL_ECHO	= 0x0001;	/* ��������ʸ���򥨥����Хå� */
// const uint_t IOCTL_CRLF	= 0x0010;	/* LF��������������CR���ղ� */
// const uint_t IOCTL_FCSND = 0x0100;	/* �������Ф��ƥե������Ԥ� */
// const uint_t IOCTL_FCANY = 0x0200;	/* �ɤΤ褦��ʸ���Ǥ������Ƴ� */
// const uint_t IOCTL_FCRCV = 0x0400;	/* �������Ф��ƥե������Ԥ� */
// ------------------------------------------+

celltype tSerialPortWrapper {
	entry sSerialPort	eSerialPort;
	entry snSerialPort	enSerialPort;
// +---  ---------------------
//  	call sSIOPort		cSIOPort;	/* �ʰ�SIO�ɥ饤�ФȤ���³ */
// 	entry siSIOCBR		eiSIOCBR;
// 	call sSemaphore  cSendSemaphore;
// 	call siSemaphore ciSendSemaphore;
// ----------------------  ---+	
    attr {
		ID   portid;
	};
};
